`ifndef SPI_UVC_TYPES_SV
`define SPI_UVC_TYPES_SV

typedef enum {
  SPI_UVC_WRITE,
  SPI_UVC_READ
} spi_uvc_cmd_e;

`endif // SPI_UVC_TYPES_SV
