`ifndef SPI_UVC_PKG_SV
`define SPI_UVC_PKG_SV

package spi_uvc_pkg;

  `include "uvm_macros.svh"
  import uvm_pkg::*;

  `include "spi_uvc_agent.sv"

endpackage : spi_uvc_pkg

`endif // SPI_UVC_PKG_SV